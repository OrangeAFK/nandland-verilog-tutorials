module example_and_gate (
    input i1, input i2,
    output and_result
);
    assign and_result = i1 & i2;

endmodule